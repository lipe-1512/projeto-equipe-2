module controlUnit (
    input clk, resert,
    
    output reg PCWrite,
    output reg PCWriteCond,
    output reg IorD,
    output reg MemWR,
    output reg IRWrite,
    output reg RegRs,
    output reg [1:0] RegDst,
    output reg RegWrite,
    output reg WrA,
    output reg WrB,
    output reg [1:0] ALUSrcA,
    output reg [1:0] ALUSrcB,
    output reg [2:0] ALUControl,
    output reg ALUOutCtrl,
    output reg EPCCtrl,
    output reg [2:0] PcSource,
    output reg [1:0] Exception,
    output reg [4:0] DataSrc,
    output reg LSControl,
    output reg SSControl,
    output reg MemDataWrite,
    output reg SEControl,
    output reg ShiftSrc,
    output reg ShiftAmt,
    output reg [2:0] ShiftControl,
    output reg MDControl,
    output reg WriteHI,
    output reg WriteLO,
    output reg div0,
    output reg resert_out,
    output reg overflow_flag,
    output reg maior_flag,
    output reg igual_flag,
    output reg menor_flag,
    output reg zero_flag
);
    
endmodule